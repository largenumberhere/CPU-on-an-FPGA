module Not(
    input in,
    output out
);
    Nand(in, 1, out);
endmodule